library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


use work.alu_pkg.all; 

entity top_alu is
generic (
  CLK_FREQ_HZ : integer := 125_000_000;
  BAUD        : integer := 115200
);
  port(
    clk            : in  std_logic;
    rst_n          : in  std_logic;
   
    btn_a_up       : in  std_logic;
    btn_a_down     : in  std_logic;
    btn_b_up       : in  std_logic;
    btn_b_down     : in  std_logic;

    -- PWM RGB
    pwm_r_o        : out std_logic;
    pwm_g_o        : out std_logic;
    pwm_b_o        : out std_logic
  );
end entity;

architecture rtl of top_alu is 
--  ----------------------------------------------------------------------------
  -- Debounced pulses
  signal a_up_p, a_dn_p, b_up_p, b_dn_p : std_logic;

  -- A/B regs 
  signal reg_a, reg_b : unsigned(7 downto 0) := (others=>'0');

  --  A/B btns
  signal btn_a_q, btn_b_q : std_logic_vector(7 downto 0);



  signal Y          : std_logic_vector(15 downto 0);

  signal duty_r, duty_g, duty_b : std_logic_vector(7 downto 0);
    
 begin


--   ----------------------------------------------------------------------------
--   -- Buttons → pulses
  db_aup : entity work.debounce_onepulse generic map(N_SAMPLES=>20000) port map(clk,rst_n,btn_a_up ,a_up_p);
  db_adn : entity work.debounce_onepulse generic map(N_SAMPLES=>20000) port map(clk,rst_n,btn_a_down,a_dn_p);
  db_bup : entity work.debounce_onepulse generic map(N_SAMPLES=>20000) port map(clk,rst_n,btn_b_up ,b_up_p);
  db_bdn : entity work.debounce_onepulse generic map(N_SAMPLES=>20000) port map(clk,rst_n,btn_b_down,b_dn_p);
  db_op : entity work.debounce_onepulse generic map(N_SAMPLES=>20000) port map(clk, rst_n, op_next, op_pulse);

  regA_btn: entity work.updown_byte port map(clk,rst_n,a_up_p,a_dn_p,btn_a_q);
  regB_btn: entity work.updown_byte port map(clk,rst_n,b_up_p,b_dn_p,btn_b_q);


  process(clk, rst_n) begin
    if rst_n='0' then
      reg_a <= (others=>'0');
      reg_b <= (others=>'0');
      op_sel <= OP_ADD;
    elsif rising_edge(clk) then
    reg_a <= unsigned(btn_a_q);
    reg_b <= unsigned(btn_b_q);
    if op_pulse='1' then
      if op_idx = "101" then     
        op_idx <= (others=>'0'); 
      else
        op_idx <= op_idx + 1;
      end if;
    end if;
    case op_idx is
      when "000" => op_sel <= OP_ADD; 
      when "001" => op_sel <= OP_SUB; 
      when "010" => op_sel <= OP_MUL; 
      when "011" => op_sel <= OP_SHL; 
      when "100" => op_sel <= OP_SHR; 
      when "101" => op_sel <= OP_SAR; 
      when others => op_sel <= OP_ADD;
    end case;
  end if;

  end process;



  duty_r <= std_logic_vector(unsigned(Y(15 downto 8)));  
  duty_g <= std_logic_vector(unsigned(Y(7 downto 0)));   
  duty_b <= std_logic_vector(unsigned(Y(7 downto 0)));        

  -- PWM  
 u_pwm_r: entity work.pwm8 port map(clk=>clk, rst_n=>rst_n, duty => duty_r , pwm => pwm_r_o);
 u_pwm_g: entity work.pwm8 port map(clk=>clk, rst_n=>rst_n, duty => duty_g , pwm => pwm_g_o);
 u_pwm_b: entity work.pwm8 port map(clk=>clk, rst_n=>rst_n, duty => duty_b , pwm => pwm_b_o);
end architecture;
