class dxi_slave_seq #(int DW=8) extends uvm_sequence #(dxi_transation#(DW));
  `uvm_object_param_utils(dxi_slave_seq#(DW))

      rand int unsigned n_items;
  constraint c_n_items { n_items inside {[50:200]}; } 


  function new(string name="dxi_slave_seq");
    super.new(name);
  endfunction

  task body();
    dxi_transation#(DW) tr;

    if (starting_phase != null)
      starting_phase.raise_objection(this);

    repeat (200) begin
      tr = dxi_transation#(DW)::type_id::create("tr");

      start_item(tr);

      if (!tr.randomize()) begin
        `uvm_fatal(get_type_name(), "Slave: tr.randomize() failed")
      end

      finish_item(tr);
    end

    if (starting_phase != null)
      starting_phase.drop_objection(this);
  endtask
endclass
