interface config_if(input logic clk);
  logic [1:0] config_select;
endinterface
