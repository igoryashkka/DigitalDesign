library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package driver_pkg is
  constant SEG_A : std_logic_vector(7 downto 0) := x"77";
  constant SEG_B : std_logic_vector(7 downto 0) := x"7C";
  constant SEG_C : std_logic_vector(7 downto 0) := x"39";
  constant SEG_D : std_logic_vector(7 downto 0) := x"3F";
  constant SEG_E : std_logic_vector(7 downto 0) := x"79";
  constant SEG_F : std_logic_vector(7 downto 0) := x"71";
  constant SEG_G : std_logic_vector(7 downto 0) := x"3D";
  constant SEG_H : std_logic_vector(7 downto 0) := x"76";
  constant SEG_J : std_logic_vector(7 downto 0) := x"1E";
  constant SEG_L : std_logic_vector(7 downto 0) := x"38";
  constant SEG_N : std_logic_vector(7 downto 0) := x"37";
  constant SEG_O : std_logic_vector(7 downto 0) := x"3F";
  constant SEG_P : std_logic_vector(7 downto 0) := x"73";
  constant SEG_S : std_logic_vector(7 downto 0) := x"6D";
  constant SEG_U : std_logic_vector(7 downto 0) := x"3E";
  constant SEG_Y : std_logic_vector(7 downto 0) := x"6E";
  constant SEG_0 : std_logic_vector(7 downto 0) := x"3F";
  constant SEG_1 : std_logic_vector(7 downto 0) := x"06";
  constant SEG_2 : std_logic_vector(7 downto 0) := x"5B";
  constant SEG_3 : std_logic_vector(7 downto 0) := x"4F";
  constant SEG_4 : std_logic_vector(7 downto 0) := x"66";
  constant SEG_5 : std_logic_vector(7 downto 0) := x"6D";
  constant SEG_6 : std_logic_vector(7 downto 0) := x"7D";
  constant SEG_7 : std_logic_vector(7 downto 0) := x"07";
  constant SEG_8 : std_logic_vector(7 downto 0) := x"7F";
  constant SEG_9 : std_logic_vector(7 downto 0) := x"6F";

end package driver_pkg;

package body driver_pkg is
end package body driver_pkg;
